
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h5e263011;
    ram_cell[       1] = 32'h0;  // 32'h15fce98f;
    ram_cell[       2] = 32'h0;  // 32'h58be6bf2;
    ram_cell[       3] = 32'h0;  // 32'haef8ed6c;
    ram_cell[       4] = 32'h0;  // 32'h0bf4bc66;
    ram_cell[       5] = 32'h0;  // 32'hd23dae33;
    ram_cell[       6] = 32'h0;  // 32'ha3762096;
    ram_cell[       7] = 32'h0;  // 32'h6dd13459;
    ram_cell[       8] = 32'h0;  // 32'hd34e39d7;
    ram_cell[       9] = 32'h0;  // 32'h4d5bc3f9;
    ram_cell[      10] = 32'h0;  // 32'h2885224f;
    ram_cell[      11] = 32'h0;  // 32'h32aa24a2;
    ram_cell[      12] = 32'h0;  // 32'ha3710f8e;
    ram_cell[      13] = 32'h0;  // 32'h0c2fc509;
    ram_cell[      14] = 32'h0;  // 32'h3675b566;
    ram_cell[      15] = 32'h0;  // 32'h26be296f;
    ram_cell[      16] = 32'h0;  // 32'hf034f6a6;
    ram_cell[      17] = 32'h0;  // 32'hef0334d4;
    ram_cell[      18] = 32'h0;  // 32'hae23d46d;
    ram_cell[      19] = 32'h0;  // 32'h7e392201;
    ram_cell[      20] = 32'h0;  // 32'h4d05c3c3;
    ram_cell[      21] = 32'h0;  // 32'hd0488cec;
    ram_cell[      22] = 32'h0;  // 32'ha734be0d;
    ram_cell[      23] = 32'h0;  // 32'h27b5b241;
    ram_cell[      24] = 32'h0;  // 32'h9a69f06c;
    ram_cell[      25] = 32'h0;  // 32'hdd56010a;
    ram_cell[      26] = 32'h0;  // 32'h1a8b5029;
    ram_cell[      27] = 32'h0;  // 32'hc50ab0d0;
    ram_cell[      28] = 32'h0;  // 32'h5b81d28b;
    ram_cell[      29] = 32'h0;  // 32'hd038c823;
    ram_cell[      30] = 32'h0;  // 32'h4cf4add0;
    ram_cell[      31] = 32'h0;  // 32'h2e2f19d7;
    ram_cell[      32] = 32'h0;  // 32'h966fe14b;
    ram_cell[      33] = 32'h0;  // 32'hb63426ba;
    ram_cell[      34] = 32'h0;  // 32'h62ea3535;
    ram_cell[      35] = 32'h0;  // 32'h0340bbd1;
    ram_cell[      36] = 32'h0;  // 32'hd1be3230;
    ram_cell[      37] = 32'h0;  // 32'hec354c77;
    ram_cell[      38] = 32'h0;  // 32'hb7eeee8a;
    ram_cell[      39] = 32'h0;  // 32'h4a5f945f;
    ram_cell[      40] = 32'h0;  // 32'hfab5e1f6;
    ram_cell[      41] = 32'h0;  // 32'hd499ac88;
    ram_cell[      42] = 32'h0;  // 32'h264d64bc;
    ram_cell[      43] = 32'h0;  // 32'h1331c782;
    ram_cell[      44] = 32'h0;  // 32'h1fe8f917;
    ram_cell[      45] = 32'h0;  // 32'ha7601a53;
    ram_cell[      46] = 32'h0;  // 32'h2bbbc698;
    ram_cell[      47] = 32'h0;  // 32'hd60904bb;
    ram_cell[      48] = 32'h0;  // 32'h1bccf3fc;
    ram_cell[      49] = 32'h0;  // 32'hfea5c3c8;
    ram_cell[      50] = 32'h0;  // 32'h1102a521;
    ram_cell[      51] = 32'h0;  // 32'hffcb0c83;
    ram_cell[      52] = 32'h0;  // 32'hc0233c41;
    ram_cell[      53] = 32'h0;  // 32'h64f921d2;
    ram_cell[      54] = 32'h0;  // 32'h9ad57759;
    ram_cell[      55] = 32'h0;  // 32'h1120b984;
    ram_cell[      56] = 32'h0;  // 32'h6e3fc592;
    ram_cell[      57] = 32'h0;  // 32'hb54d64f7;
    ram_cell[      58] = 32'h0;  // 32'h27f9ce42;
    ram_cell[      59] = 32'h0;  // 32'hd97b76ef;
    ram_cell[      60] = 32'h0;  // 32'h3cab69d7;
    ram_cell[      61] = 32'h0;  // 32'hc319fefd;
    ram_cell[      62] = 32'h0;  // 32'hcfa3140a;
    ram_cell[      63] = 32'h0;  // 32'hbbbb7fe6;
    ram_cell[      64] = 32'h0;  // 32'h12b8b59d;
    ram_cell[      65] = 32'h0;  // 32'hc1d5c7ec;
    ram_cell[      66] = 32'h0;  // 32'h36ed5af8;
    ram_cell[      67] = 32'h0;  // 32'hdb101abc;
    ram_cell[      68] = 32'h0;  // 32'h05f13329;
    ram_cell[      69] = 32'h0;  // 32'h55330ea3;
    ram_cell[      70] = 32'h0;  // 32'h78a9559a;
    ram_cell[      71] = 32'h0;  // 32'h0f567021;
    ram_cell[      72] = 32'h0;  // 32'h983284b9;
    ram_cell[      73] = 32'h0;  // 32'h993542e3;
    ram_cell[      74] = 32'h0;  // 32'hb88d2456;
    ram_cell[      75] = 32'h0;  // 32'heeb41c86;
    ram_cell[      76] = 32'h0;  // 32'hb64f0e52;
    ram_cell[      77] = 32'h0;  // 32'h525d4401;
    ram_cell[      78] = 32'h0;  // 32'h6ab7ef35;
    ram_cell[      79] = 32'h0;  // 32'h44906c87;
    ram_cell[      80] = 32'h0;  // 32'h76ef4a4f;
    ram_cell[      81] = 32'h0;  // 32'h124a475b;
    ram_cell[      82] = 32'h0;  // 32'h5640ae07;
    ram_cell[      83] = 32'h0;  // 32'ha12dd808;
    ram_cell[      84] = 32'h0;  // 32'h3dbb39fe;
    ram_cell[      85] = 32'h0;  // 32'hd7f75823;
    ram_cell[      86] = 32'h0;  // 32'h0ff48039;
    ram_cell[      87] = 32'h0;  // 32'hb83e2115;
    ram_cell[      88] = 32'h0;  // 32'he660fb00;
    ram_cell[      89] = 32'h0;  // 32'h292e56bb;
    ram_cell[      90] = 32'h0;  // 32'hd93da5a8;
    ram_cell[      91] = 32'h0;  // 32'h67419df3;
    ram_cell[      92] = 32'h0;  // 32'h029afbf8;
    ram_cell[      93] = 32'h0;  // 32'h4d89c59f;
    ram_cell[      94] = 32'h0;  // 32'h7539afdd;
    ram_cell[      95] = 32'h0;  // 32'hea167b4e;
    ram_cell[      96] = 32'h0;  // 32'h463d7136;
    ram_cell[      97] = 32'h0;  // 32'ha1829af5;
    ram_cell[      98] = 32'h0;  // 32'h06d7e1d5;
    ram_cell[      99] = 32'h0;  // 32'h5e1512a8;
    ram_cell[     100] = 32'h0;  // 32'h0fbb539b;
    ram_cell[     101] = 32'h0;  // 32'h0db90367;
    ram_cell[     102] = 32'h0;  // 32'h75a97492;
    ram_cell[     103] = 32'h0;  // 32'h0afdbf8d;
    ram_cell[     104] = 32'h0;  // 32'he2a5420c;
    ram_cell[     105] = 32'h0;  // 32'h0d4ed830;
    ram_cell[     106] = 32'h0;  // 32'hd5f92c46;
    ram_cell[     107] = 32'h0;  // 32'hc9d233c9;
    ram_cell[     108] = 32'h0;  // 32'hf2d36368;
    ram_cell[     109] = 32'h0;  // 32'h37d5a5de;
    ram_cell[     110] = 32'h0;  // 32'hdf88ada7;
    ram_cell[     111] = 32'h0;  // 32'h45c48caa;
    ram_cell[     112] = 32'h0;  // 32'h8af776e1;
    ram_cell[     113] = 32'h0;  // 32'h8f0790ac;
    ram_cell[     114] = 32'h0;  // 32'h285a3317;
    ram_cell[     115] = 32'h0;  // 32'hfdd77d4b;
    ram_cell[     116] = 32'h0;  // 32'h4d0f7c7a;
    ram_cell[     117] = 32'h0;  // 32'hc8e28142;
    ram_cell[     118] = 32'h0;  // 32'hcb6dc468;
    ram_cell[     119] = 32'h0;  // 32'hdbd31181;
    ram_cell[     120] = 32'h0;  // 32'h94645f21;
    ram_cell[     121] = 32'h0;  // 32'h93ae59b9;
    ram_cell[     122] = 32'h0;  // 32'hdb509377;
    ram_cell[     123] = 32'h0;  // 32'hfdda9489;
    ram_cell[     124] = 32'h0;  // 32'h0f0f73e2;
    ram_cell[     125] = 32'h0;  // 32'hb89e3093;
    ram_cell[     126] = 32'h0;  // 32'h30a21534;
    ram_cell[     127] = 32'h0;  // 32'he825dd6f;
    ram_cell[     128] = 32'h0;  // 32'h9d3d381f;
    ram_cell[     129] = 32'h0;  // 32'h021118af;
    ram_cell[     130] = 32'h0;  // 32'h7a8e0788;
    ram_cell[     131] = 32'h0;  // 32'h02551262;
    ram_cell[     132] = 32'h0;  // 32'hecfa861a;
    ram_cell[     133] = 32'h0;  // 32'he1576071;
    ram_cell[     134] = 32'h0;  // 32'h67cde764;
    ram_cell[     135] = 32'h0;  // 32'he1428ac4;
    ram_cell[     136] = 32'h0;  // 32'h83be28c8;
    ram_cell[     137] = 32'h0;  // 32'h3c985c6d;
    ram_cell[     138] = 32'h0;  // 32'h3634d632;
    ram_cell[     139] = 32'h0;  // 32'hb31c5c5d;
    ram_cell[     140] = 32'h0;  // 32'h46445a56;
    ram_cell[     141] = 32'h0;  // 32'h934ee19e;
    ram_cell[     142] = 32'h0;  // 32'h478e1726;
    ram_cell[     143] = 32'h0;  // 32'hebcb51de;
    ram_cell[     144] = 32'h0;  // 32'h43a5690a;
    ram_cell[     145] = 32'h0;  // 32'he9d829cb;
    ram_cell[     146] = 32'h0;  // 32'h2e4155b0;
    ram_cell[     147] = 32'h0;  // 32'hcc9beeb9;
    ram_cell[     148] = 32'h0;  // 32'hb3ab7fae;
    ram_cell[     149] = 32'h0;  // 32'h06ede333;
    ram_cell[     150] = 32'h0;  // 32'h004f93bb;
    ram_cell[     151] = 32'h0;  // 32'h9480d922;
    ram_cell[     152] = 32'h0;  // 32'h6cad5a6d;
    ram_cell[     153] = 32'h0;  // 32'h6804e83e;
    ram_cell[     154] = 32'h0;  // 32'hd350691a;
    ram_cell[     155] = 32'h0;  // 32'h10f9af40;
    ram_cell[     156] = 32'h0;  // 32'ha1b8a9d3;
    ram_cell[     157] = 32'h0;  // 32'hcaf53a9e;
    ram_cell[     158] = 32'h0;  // 32'ha8aa677d;
    ram_cell[     159] = 32'h0;  // 32'h1e987425;
    ram_cell[     160] = 32'h0;  // 32'h8c564731;
    ram_cell[     161] = 32'h0;  // 32'h7c7a88be;
    ram_cell[     162] = 32'h0;  // 32'hb9d1f512;
    ram_cell[     163] = 32'h0;  // 32'h6d8a75be;
    ram_cell[     164] = 32'h0;  // 32'h1721c23f;
    ram_cell[     165] = 32'h0;  // 32'he2857a3e;
    ram_cell[     166] = 32'h0;  // 32'h0afeefe6;
    ram_cell[     167] = 32'h0;  // 32'h63ecf667;
    ram_cell[     168] = 32'h0;  // 32'h54b0e579;
    ram_cell[     169] = 32'h0;  // 32'hb40afc42;
    ram_cell[     170] = 32'h0;  // 32'hbdc325c0;
    ram_cell[     171] = 32'h0;  // 32'h695b6efb;
    ram_cell[     172] = 32'h0;  // 32'hc7869b4c;
    ram_cell[     173] = 32'h0;  // 32'h707630fc;
    ram_cell[     174] = 32'h0;  // 32'h28f0492d;
    ram_cell[     175] = 32'h0;  // 32'h9ca61ece;
    ram_cell[     176] = 32'h0;  // 32'hefcc31eb;
    ram_cell[     177] = 32'h0;  // 32'h780aaa7c;
    ram_cell[     178] = 32'h0;  // 32'h68f06de0;
    ram_cell[     179] = 32'h0;  // 32'hf8d6235b;
    ram_cell[     180] = 32'h0;  // 32'h972e22a0;
    ram_cell[     181] = 32'h0;  // 32'h76690580;
    ram_cell[     182] = 32'h0;  // 32'h40369823;
    ram_cell[     183] = 32'h0;  // 32'h29cab230;
    ram_cell[     184] = 32'h0;  // 32'h42f64f87;
    ram_cell[     185] = 32'h0;  // 32'h3d942255;
    ram_cell[     186] = 32'h0;  // 32'hc1e29ff0;
    ram_cell[     187] = 32'h0;  // 32'hbf5e2079;
    ram_cell[     188] = 32'h0;  // 32'h6bbe5fe4;
    ram_cell[     189] = 32'h0;  // 32'hfbff9849;
    ram_cell[     190] = 32'h0;  // 32'h13b110be;
    ram_cell[     191] = 32'h0;  // 32'hb5ab4d98;
    ram_cell[     192] = 32'h0;  // 32'h0e27fe8b;
    ram_cell[     193] = 32'h0;  // 32'h9b344958;
    ram_cell[     194] = 32'h0;  // 32'h9911164d;
    ram_cell[     195] = 32'h0;  // 32'h98a38abc;
    ram_cell[     196] = 32'h0;  // 32'h19dc6459;
    ram_cell[     197] = 32'h0;  // 32'h751ff77d;
    ram_cell[     198] = 32'h0;  // 32'h3a7a06c8;
    ram_cell[     199] = 32'h0;  // 32'h28d3795d;
    ram_cell[     200] = 32'h0;  // 32'ha651efcc;
    ram_cell[     201] = 32'h0;  // 32'h2d6a91cc;
    ram_cell[     202] = 32'h0;  // 32'h153009a1;
    ram_cell[     203] = 32'h0;  // 32'hff56c195;
    ram_cell[     204] = 32'h0;  // 32'h00a8eadb;
    ram_cell[     205] = 32'h0;  // 32'h2f9704e9;
    ram_cell[     206] = 32'h0;  // 32'h9cdb671b;
    ram_cell[     207] = 32'h0;  // 32'h5beb50ad;
    ram_cell[     208] = 32'h0;  // 32'hdd7797ec;
    ram_cell[     209] = 32'h0;  // 32'h37ffad8f;
    ram_cell[     210] = 32'h0;  // 32'hb660f0f5;
    ram_cell[     211] = 32'h0;  // 32'he039f476;
    ram_cell[     212] = 32'h0;  // 32'hce23860c;
    ram_cell[     213] = 32'h0;  // 32'h0780233d;
    ram_cell[     214] = 32'h0;  // 32'hf469619b;
    ram_cell[     215] = 32'h0;  // 32'h5e738966;
    ram_cell[     216] = 32'h0;  // 32'hb5a24b72;
    ram_cell[     217] = 32'h0;  // 32'hcc77f95a;
    ram_cell[     218] = 32'h0;  // 32'h273ceb20;
    ram_cell[     219] = 32'h0;  // 32'he202f0ea;
    ram_cell[     220] = 32'h0;  // 32'h2718aeab;
    ram_cell[     221] = 32'h0;  // 32'h6e786234;
    ram_cell[     222] = 32'h0;  // 32'h6020d6c9;
    ram_cell[     223] = 32'h0;  // 32'h74337cbb;
    ram_cell[     224] = 32'h0;  // 32'h9ca12e7a;
    ram_cell[     225] = 32'h0;  // 32'h67a5f6b9;
    ram_cell[     226] = 32'h0;  // 32'h14d7c7d7;
    ram_cell[     227] = 32'h0;  // 32'h20b55c36;
    ram_cell[     228] = 32'h0;  // 32'h089ac54d;
    ram_cell[     229] = 32'h0;  // 32'hde11a5a8;
    ram_cell[     230] = 32'h0;  // 32'h4618f161;
    ram_cell[     231] = 32'h0;  // 32'ha925113a;
    ram_cell[     232] = 32'h0;  // 32'hd1c941c0;
    ram_cell[     233] = 32'h0;  // 32'h15d32309;
    ram_cell[     234] = 32'h0;  // 32'hb4331de6;
    ram_cell[     235] = 32'h0;  // 32'h77b8b0b4;
    ram_cell[     236] = 32'h0;  // 32'h0154f861;
    ram_cell[     237] = 32'h0;  // 32'hc5d6b473;
    ram_cell[     238] = 32'h0;  // 32'hf8b38990;
    ram_cell[     239] = 32'h0;  // 32'h22cb6344;
    ram_cell[     240] = 32'h0;  // 32'h0e9ea05e;
    ram_cell[     241] = 32'h0;  // 32'hc48024f1;
    ram_cell[     242] = 32'h0;  // 32'h2bbe8cd9;
    ram_cell[     243] = 32'h0;  // 32'h10d4a802;
    ram_cell[     244] = 32'h0;  // 32'hf875ded5;
    ram_cell[     245] = 32'h0;  // 32'hf337b79d;
    ram_cell[     246] = 32'h0;  // 32'h38f7c12c;
    ram_cell[     247] = 32'h0;  // 32'h6dfc9188;
    ram_cell[     248] = 32'h0;  // 32'h46ce975e;
    ram_cell[     249] = 32'h0;  // 32'hd4760320;
    ram_cell[     250] = 32'h0;  // 32'h4fb496f5;
    ram_cell[     251] = 32'h0;  // 32'h11190396;
    ram_cell[     252] = 32'h0;  // 32'hd9eb047a;
    ram_cell[     253] = 32'h0;  // 32'h1cf4c438;
    ram_cell[     254] = 32'h0;  // 32'hb47cff31;
    ram_cell[     255] = 32'h0;  // 32'hfd50ce7e;
    // src matrix A
    ram_cell[     256] = 32'hd9a56d9a;
    ram_cell[     257] = 32'hfce2eb41;
    ram_cell[     258] = 32'hc49e6482;
    ram_cell[     259] = 32'h569d1ed5;
    ram_cell[     260] = 32'h0e4ce5fa;
    ram_cell[     261] = 32'h8c628f2c;
    ram_cell[     262] = 32'h6041b57e;
    ram_cell[     263] = 32'h57c1c6d2;
    ram_cell[     264] = 32'hc207ebab;
    ram_cell[     265] = 32'hf8380c4e;
    ram_cell[     266] = 32'h86fa2489;
    ram_cell[     267] = 32'h0fa53bae;
    ram_cell[     268] = 32'hf8bdc73c;
    ram_cell[     269] = 32'ha80fe0f5;
    ram_cell[     270] = 32'ha301c1ef;
    ram_cell[     271] = 32'h5f92f944;
    ram_cell[     272] = 32'h6284ea99;
    ram_cell[     273] = 32'h2388f356;
    ram_cell[     274] = 32'hae25ae1f;
    ram_cell[     275] = 32'h740894fb;
    ram_cell[     276] = 32'h44b03598;
    ram_cell[     277] = 32'h97455849;
    ram_cell[     278] = 32'h2ab39f58;
    ram_cell[     279] = 32'h682871a5;
    ram_cell[     280] = 32'hc4299358;
    ram_cell[     281] = 32'h128cee7e;
    ram_cell[     282] = 32'h3c15f682;
    ram_cell[     283] = 32'hd92a1574;
    ram_cell[     284] = 32'h7d381a15;
    ram_cell[     285] = 32'he95d8b56;
    ram_cell[     286] = 32'hd9e61301;
    ram_cell[     287] = 32'hd7bde109;
    ram_cell[     288] = 32'hd099433f;
    ram_cell[     289] = 32'h80763f47;
    ram_cell[     290] = 32'h546955d8;
    ram_cell[     291] = 32'hc7fd2210;
    ram_cell[     292] = 32'h3184ed18;
    ram_cell[     293] = 32'hc48bb8a2;
    ram_cell[     294] = 32'hb086768a;
    ram_cell[     295] = 32'h0457a5f6;
    ram_cell[     296] = 32'he89bfc16;
    ram_cell[     297] = 32'hb9ef7cee;
    ram_cell[     298] = 32'hc390e96d;
    ram_cell[     299] = 32'h57822ebb;
    ram_cell[     300] = 32'h92242316;
    ram_cell[     301] = 32'hb7bed005;
    ram_cell[     302] = 32'h2803e043;
    ram_cell[     303] = 32'h9b80e8e5;
    ram_cell[     304] = 32'h08bbb22c;
    ram_cell[     305] = 32'hb1411b36;
    ram_cell[     306] = 32'h5bd157c0;
    ram_cell[     307] = 32'hf624f6ee;
    ram_cell[     308] = 32'h61bfdaee;
    ram_cell[     309] = 32'h2b53490f;
    ram_cell[     310] = 32'hc6dc9380;
    ram_cell[     311] = 32'h1fe8f1ef;
    ram_cell[     312] = 32'h1d8883d3;
    ram_cell[     313] = 32'h31c55a8d;
    ram_cell[     314] = 32'h266a630b;
    ram_cell[     315] = 32'hc9692036;
    ram_cell[     316] = 32'h0430bd60;
    ram_cell[     317] = 32'h7353fcc4;
    ram_cell[     318] = 32'h18c602e0;
    ram_cell[     319] = 32'h4cc50939;
    ram_cell[     320] = 32'hf6576ba1;
    ram_cell[     321] = 32'h18e4567c;
    ram_cell[     322] = 32'h0e201ac6;
    ram_cell[     323] = 32'hde3edc47;
    ram_cell[     324] = 32'h356e26c5;
    ram_cell[     325] = 32'h3f59869b;
    ram_cell[     326] = 32'h399a96b6;
    ram_cell[     327] = 32'h3b06a740;
    ram_cell[     328] = 32'hae8fa18f;
    ram_cell[     329] = 32'h0b9bf8cc;
    ram_cell[     330] = 32'hf64f2d9e;
    ram_cell[     331] = 32'h0bcc224a;
    ram_cell[     332] = 32'h78174974;
    ram_cell[     333] = 32'h43da7205;
    ram_cell[     334] = 32'h88db0ee4;
    ram_cell[     335] = 32'h51011db3;
    ram_cell[     336] = 32'h71ee756e;
    ram_cell[     337] = 32'h86b0ed22;
    ram_cell[     338] = 32'hb553ef5a;
    ram_cell[     339] = 32'h605075df;
    ram_cell[     340] = 32'h9051a332;
    ram_cell[     341] = 32'h679a72f6;
    ram_cell[     342] = 32'h8aa73368;
    ram_cell[     343] = 32'hfbab2094;
    ram_cell[     344] = 32'h2430e927;
    ram_cell[     345] = 32'h845f6b06;
    ram_cell[     346] = 32'h3558c73b;
    ram_cell[     347] = 32'hfbb0b533;
    ram_cell[     348] = 32'hb2915f4f;
    ram_cell[     349] = 32'hef7a4425;
    ram_cell[     350] = 32'hee9e1846;
    ram_cell[     351] = 32'hef95d744;
    ram_cell[     352] = 32'h858c8ac7;
    ram_cell[     353] = 32'h6951fd2c;
    ram_cell[     354] = 32'hf19da35a;
    ram_cell[     355] = 32'h1d8e54f1;
    ram_cell[     356] = 32'h14accbba;
    ram_cell[     357] = 32'h41cec870;
    ram_cell[     358] = 32'hccdfa361;
    ram_cell[     359] = 32'h64a8fc07;
    ram_cell[     360] = 32'h0d9d8252;
    ram_cell[     361] = 32'hb71dfb99;
    ram_cell[     362] = 32'h32452bc0;
    ram_cell[     363] = 32'hd2bcffe3;
    ram_cell[     364] = 32'h28813efb;
    ram_cell[     365] = 32'h7a225eb6;
    ram_cell[     366] = 32'h00c1ca36;
    ram_cell[     367] = 32'hcd6bdf8f;
    ram_cell[     368] = 32'h441bd417;
    ram_cell[     369] = 32'h22ac9f7a;
    ram_cell[     370] = 32'hf00865fa;
    ram_cell[     371] = 32'h3c1e3b78;
    ram_cell[     372] = 32'hc6fa0a21;
    ram_cell[     373] = 32'h07966661;
    ram_cell[     374] = 32'h368565cc;
    ram_cell[     375] = 32'h27a345e4;
    ram_cell[     376] = 32'h7afa2671;
    ram_cell[     377] = 32'h4c72d9f8;
    ram_cell[     378] = 32'hc1d4a8f3;
    ram_cell[     379] = 32'h11bd290f;
    ram_cell[     380] = 32'h1bcaf926;
    ram_cell[     381] = 32'h1d7f90f6;
    ram_cell[     382] = 32'h23ed2676;
    ram_cell[     383] = 32'h12ea2597;
    ram_cell[     384] = 32'hec395b20;
    ram_cell[     385] = 32'ha96ecaad;
    ram_cell[     386] = 32'habb112c6;
    ram_cell[     387] = 32'h660a584e;
    ram_cell[     388] = 32'hf2eadd8a;
    ram_cell[     389] = 32'h0af5592d;
    ram_cell[     390] = 32'h2f170391;
    ram_cell[     391] = 32'ha8a8a5f9;
    ram_cell[     392] = 32'h759b8557;
    ram_cell[     393] = 32'hfb0a9f47;
    ram_cell[     394] = 32'h80659967;
    ram_cell[     395] = 32'h10e46e86;
    ram_cell[     396] = 32'h9739b097;
    ram_cell[     397] = 32'h5c443f41;
    ram_cell[     398] = 32'h5e20b003;
    ram_cell[     399] = 32'h338a61a5;
    ram_cell[     400] = 32'hee758d32;
    ram_cell[     401] = 32'h219dbc9d;
    ram_cell[     402] = 32'h9c839774;
    ram_cell[     403] = 32'h74c5622c;
    ram_cell[     404] = 32'h4dd06cdb;
    ram_cell[     405] = 32'ha6d69feb;
    ram_cell[     406] = 32'he8e874f2;
    ram_cell[     407] = 32'h062e0496;
    ram_cell[     408] = 32'hd376aee7;
    ram_cell[     409] = 32'heb8acf1b;
    ram_cell[     410] = 32'h755309dc;
    ram_cell[     411] = 32'h41c58463;
    ram_cell[     412] = 32'h06221934;
    ram_cell[     413] = 32'h6b81cadd;
    ram_cell[     414] = 32'hf2bb1aec;
    ram_cell[     415] = 32'h093fec62;
    ram_cell[     416] = 32'h46f8d094;
    ram_cell[     417] = 32'h3b927ec0;
    ram_cell[     418] = 32'h73faa281;
    ram_cell[     419] = 32'h34e25a0d;
    ram_cell[     420] = 32'h32b19754;
    ram_cell[     421] = 32'hd85f0fd9;
    ram_cell[     422] = 32'h57b7d4c7;
    ram_cell[     423] = 32'he3d0c6d3;
    ram_cell[     424] = 32'h80acada1;
    ram_cell[     425] = 32'h5b6b8d79;
    ram_cell[     426] = 32'ha04df99c;
    ram_cell[     427] = 32'h51f38afa;
    ram_cell[     428] = 32'h8ad991fd;
    ram_cell[     429] = 32'hc7be568c;
    ram_cell[     430] = 32'hcd7feb11;
    ram_cell[     431] = 32'h6795f4a7;
    ram_cell[     432] = 32'hd2f62724;
    ram_cell[     433] = 32'h5ecbe649;
    ram_cell[     434] = 32'hae73ec26;
    ram_cell[     435] = 32'hee37a142;
    ram_cell[     436] = 32'h899beebb;
    ram_cell[     437] = 32'h24f1a5ee;
    ram_cell[     438] = 32'hba01e7c4;
    ram_cell[     439] = 32'hf8af1eb2;
    ram_cell[     440] = 32'hf982240c;
    ram_cell[     441] = 32'h4ee91fd0;
    ram_cell[     442] = 32'hb3d54701;
    ram_cell[     443] = 32'h6fbffd63;
    ram_cell[     444] = 32'hdc17471f;
    ram_cell[     445] = 32'hfbc745bd;
    ram_cell[     446] = 32'h58816987;
    ram_cell[     447] = 32'hf2dc7785;
    ram_cell[     448] = 32'haa9563d7;
    ram_cell[     449] = 32'h14adb01c;
    ram_cell[     450] = 32'h187443a5;
    ram_cell[     451] = 32'h4eac8c5e;
    ram_cell[     452] = 32'h73158e75;
    ram_cell[     453] = 32'h9426b883;
    ram_cell[     454] = 32'h3e13e6a7;
    ram_cell[     455] = 32'h089394df;
    ram_cell[     456] = 32'hae8e8f1e;
    ram_cell[     457] = 32'h4af2eeda;
    ram_cell[     458] = 32'h79cf5a19;
    ram_cell[     459] = 32'hbb6c500a;
    ram_cell[     460] = 32'h368558d8;
    ram_cell[     461] = 32'h52f0124a;
    ram_cell[     462] = 32'hbaa44514;
    ram_cell[     463] = 32'h225deb23;
    ram_cell[     464] = 32'h745cb1bd;
    ram_cell[     465] = 32'hc72abfbd;
    ram_cell[     466] = 32'h909e4653;
    ram_cell[     467] = 32'hc237597e;
    ram_cell[     468] = 32'h8a3e57f5;
    ram_cell[     469] = 32'hd6be96c9;
    ram_cell[     470] = 32'h521dd155;
    ram_cell[     471] = 32'h4a04af09;
    ram_cell[     472] = 32'h6a958e6c;
    ram_cell[     473] = 32'h68882b0e;
    ram_cell[     474] = 32'hd82a079f;
    ram_cell[     475] = 32'h74c70eac;
    ram_cell[     476] = 32'hd3215102;
    ram_cell[     477] = 32'h64215384;
    ram_cell[     478] = 32'h17c8b738;
    ram_cell[     479] = 32'h9df20e1c;
    ram_cell[     480] = 32'h03afaf55;
    ram_cell[     481] = 32'h9007a54e;
    ram_cell[     482] = 32'h99426b4d;
    ram_cell[     483] = 32'hc03a63c0;
    ram_cell[     484] = 32'hae29ac34;
    ram_cell[     485] = 32'hc75467f7;
    ram_cell[     486] = 32'he3556271;
    ram_cell[     487] = 32'h8e9ea16c;
    ram_cell[     488] = 32'h42ed422f;
    ram_cell[     489] = 32'ha5a68fab;
    ram_cell[     490] = 32'h87d4b630;
    ram_cell[     491] = 32'hd7acdcc1;
    ram_cell[     492] = 32'had9c260a;
    ram_cell[     493] = 32'h9af8f3cb;
    ram_cell[     494] = 32'h570ff7f4;
    ram_cell[     495] = 32'ha602ef00;
    ram_cell[     496] = 32'h1a30920b;
    ram_cell[     497] = 32'h9694cbae;
    ram_cell[     498] = 32'h4614d649;
    ram_cell[     499] = 32'hd0e0cef3;
    ram_cell[     500] = 32'h07a24bac;
    ram_cell[     501] = 32'h1a6e808c;
    ram_cell[     502] = 32'h48422fb5;
    ram_cell[     503] = 32'h726327b5;
    ram_cell[     504] = 32'h597967f8;
    ram_cell[     505] = 32'h400e8da2;
    ram_cell[     506] = 32'h86e1caf2;
    ram_cell[     507] = 32'h414aa1ac;
    ram_cell[     508] = 32'h8c44076c;
    ram_cell[     509] = 32'heea59662;
    ram_cell[     510] = 32'h0a125980;
    ram_cell[     511] = 32'hbcecd253;
    // src matrix B
    ram_cell[     512] = 32'h006e552a;
    ram_cell[     513] = 32'h6006bbd2;
    ram_cell[     514] = 32'h252c1eb8;
    ram_cell[     515] = 32'h8ed8be6d;
    ram_cell[     516] = 32'h73ef322b;
    ram_cell[     517] = 32'h0a030c2e;
    ram_cell[     518] = 32'h89c640b3;
    ram_cell[     519] = 32'h1eeb9f98;
    ram_cell[     520] = 32'h93f309e0;
    ram_cell[     521] = 32'h68f40906;
    ram_cell[     522] = 32'h8c787439;
    ram_cell[     523] = 32'hae6928f9;
    ram_cell[     524] = 32'h64c6fac9;
    ram_cell[     525] = 32'h9b6baacd;
    ram_cell[     526] = 32'he655c37a;
    ram_cell[     527] = 32'hc71c06a5;
    ram_cell[     528] = 32'hc270a00b;
    ram_cell[     529] = 32'h3b641378;
    ram_cell[     530] = 32'h3f19e000;
    ram_cell[     531] = 32'he9431af1;
    ram_cell[     532] = 32'h47d74f7d;
    ram_cell[     533] = 32'h7089c5b9;
    ram_cell[     534] = 32'hcb33aefc;
    ram_cell[     535] = 32'h8499edb0;
    ram_cell[     536] = 32'h06768286;
    ram_cell[     537] = 32'h21e11625;
    ram_cell[     538] = 32'hfd2fd74a;
    ram_cell[     539] = 32'hbed2e209;
    ram_cell[     540] = 32'h6d09fc13;
    ram_cell[     541] = 32'h280b4c76;
    ram_cell[     542] = 32'hb98dd879;
    ram_cell[     543] = 32'hc8c4d116;
    ram_cell[     544] = 32'h5553a074;
    ram_cell[     545] = 32'hafdd30d8;
    ram_cell[     546] = 32'h80e4c4a8;
    ram_cell[     547] = 32'h9a9df4fe;
    ram_cell[     548] = 32'hb634b193;
    ram_cell[     549] = 32'h39b6a164;
    ram_cell[     550] = 32'h5aa6de3c;
    ram_cell[     551] = 32'hae63aabf;
    ram_cell[     552] = 32'h6f0fff3b;
    ram_cell[     553] = 32'hf3368b21;
    ram_cell[     554] = 32'h748b142f;
    ram_cell[     555] = 32'h8b9a027c;
    ram_cell[     556] = 32'hf6a8ef69;
    ram_cell[     557] = 32'hcbec25e2;
    ram_cell[     558] = 32'hdc7f650e;
    ram_cell[     559] = 32'hffb3275b;
    ram_cell[     560] = 32'hf731a9da;
    ram_cell[     561] = 32'h2dd82f80;
    ram_cell[     562] = 32'hf0b96b42;
    ram_cell[     563] = 32'h7944c5bd;
    ram_cell[     564] = 32'hdd52a5ea;
    ram_cell[     565] = 32'hce03ca32;
    ram_cell[     566] = 32'hf84d8073;
    ram_cell[     567] = 32'hb494c4b3;
    ram_cell[     568] = 32'h7288256e;
    ram_cell[     569] = 32'h0a49c56f;
    ram_cell[     570] = 32'h8c1177a6;
    ram_cell[     571] = 32'h0455ef2a;
    ram_cell[     572] = 32'h363c3eaf;
    ram_cell[     573] = 32'h043b5515;
    ram_cell[     574] = 32'hd2a610a4;
    ram_cell[     575] = 32'h5bee7181;
    ram_cell[     576] = 32'h9d7eb67e;
    ram_cell[     577] = 32'h39aab36e;
    ram_cell[     578] = 32'hb1301fff;
    ram_cell[     579] = 32'hc752ff92;
    ram_cell[     580] = 32'hfe265a0d;
    ram_cell[     581] = 32'h6fd745c5;
    ram_cell[     582] = 32'ha4e093b2;
    ram_cell[     583] = 32'h1ec29bce;
    ram_cell[     584] = 32'hab9b90b8;
    ram_cell[     585] = 32'h3fa86c40;
    ram_cell[     586] = 32'h848708c3;
    ram_cell[     587] = 32'h69826e5b;
    ram_cell[     588] = 32'h52830a00;
    ram_cell[     589] = 32'he200286d;
    ram_cell[     590] = 32'h8766a846;
    ram_cell[     591] = 32'hfa4a46a7;
    ram_cell[     592] = 32'h4b477ff9;
    ram_cell[     593] = 32'hbefcef30;
    ram_cell[     594] = 32'h4070bee8;
    ram_cell[     595] = 32'h015bb547;
    ram_cell[     596] = 32'h09e8f462;
    ram_cell[     597] = 32'h2da1b628;
    ram_cell[     598] = 32'h05c2d40f;
    ram_cell[     599] = 32'h19c85994;
    ram_cell[     600] = 32'he2eea501;
    ram_cell[     601] = 32'h94557555;
    ram_cell[     602] = 32'h2d4bdcdc;
    ram_cell[     603] = 32'h6a34bfc3;
    ram_cell[     604] = 32'h8ebf4f43;
    ram_cell[     605] = 32'h0f22583c;
    ram_cell[     606] = 32'h454eb354;
    ram_cell[     607] = 32'h7b0af1dd;
    ram_cell[     608] = 32'he0a6df39;
    ram_cell[     609] = 32'h9ed95554;
    ram_cell[     610] = 32'hbd63c140;
    ram_cell[     611] = 32'h83fbbab9;
    ram_cell[     612] = 32'hdd773a27;
    ram_cell[     613] = 32'h8c818627;
    ram_cell[     614] = 32'he3b368ef;
    ram_cell[     615] = 32'h8bcd8bdd;
    ram_cell[     616] = 32'h18280abc;
    ram_cell[     617] = 32'hb55a5117;
    ram_cell[     618] = 32'h505677d1;
    ram_cell[     619] = 32'h0273d615;
    ram_cell[     620] = 32'h97af0349;
    ram_cell[     621] = 32'h1c0c0c43;
    ram_cell[     622] = 32'hd31f7c7c;
    ram_cell[     623] = 32'hcd25108a;
    ram_cell[     624] = 32'h39184845;
    ram_cell[     625] = 32'h647ddb80;
    ram_cell[     626] = 32'h91e431ab;
    ram_cell[     627] = 32'ha0d64bd0;
    ram_cell[     628] = 32'hf3fcd3b2;
    ram_cell[     629] = 32'h81a31f43;
    ram_cell[     630] = 32'hd9370884;
    ram_cell[     631] = 32'h8b42e1b2;
    ram_cell[     632] = 32'hae7e6d43;
    ram_cell[     633] = 32'h2d835e0c;
    ram_cell[     634] = 32'h11ccf245;
    ram_cell[     635] = 32'h4e410a88;
    ram_cell[     636] = 32'hd765f6c3;
    ram_cell[     637] = 32'h624f22ba;
    ram_cell[     638] = 32'h8ce1684a;
    ram_cell[     639] = 32'h838bb5d5;
    ram_cell[     640] = 32'haa29a6e9;
    ram_cell[     641] = 32'h455c51e9;
    ram_cell[     642] = 32'h4053f436;
    ram_cell[     643] = 32'h43d76d60;
    ram_cell[     644] = 32'hcf916405;
    ram_cell[     645] = 32'h5c352c32;
    ram_cell[     646] = 32'h6751437b;
    ram_cell[     647] = 32'h779db12e;
    ram_cell[     648] = 32'h8b0c85d7;
    ram_cell[     649] = 32'h09c90264;
    ram_cell[     650] = 32'h3dc1ab89;
    ram_cell[     651] = 32'h3f4d46db;
    ram_cell[     652] = 32'h79dcc1cc;
    ram_cell[     653] = 32'h2597091b;
    ram_cell[     654] = 32'h301b6c10;
    ram_cell[     655] = 32'h9f75a103;
    ram_cell[     656] = 32'h3d06e101;
    ram_cell[     657] = 32'h1298d4bb;
    ram_cell[     658] = 32'h75ad4779;
    ram_cell[     659] = 32'hd3ed2f9f;
    ram_cell[     660] = 32'hca2a9125;
    ram_cell[     661] = 32'ha340fe45;
    ram_cell[     662] = 32'h1d4c5e14;
    ram_cell[     663] = 32'hf9574c6d;
    ram_cell[     664] = 32'h4cf84fb4;
    ram_cell[     665] = 32'h80c7339b;
    ram_cell[     666] = 32'hf405a9cc;
    ram_cell[     667] = 32'h9959ed90;
    ram_cell[     668] = 32'h951c795b;
    ram_cell[     669] = 32'h8188d8d6;
    ram_cell[     670] = 32'he2cf8935;
    ram_cell[     671] = 32'h7fa67c47;
    ram_cell[     672] = 32'hefa74fa4;
    ram_cell[     673] = 32'hae3dcbd1;
    ram_cell[     674] = 32'hf3b148b9;
    ram_cell[     675] = 32'hb919ffa4;
    ram_cell[     676] = 32'h9881564d;
    ram_cell[     677] = 32'hb498a0f5;
    ram_cell[     678] = 32'h1fce0c96;
    ram_cell[     679] = 32'h10b8911e;
    ram_cell[     680] = 32'hf20ced07;
    ram_cell[     681] = 32'hbfdb7a84;
    ram_cell[     682] = 32'hf23df569;
    ram_cell[     683] = 32'ha8edbfdf;
    ram_cell[     684] = 32'haca38271;
    ram_cell[     685] = 32'hb9abcbbb;
    ram_cell[     686] = 32'hbb9aa86e;
    ram_cell[     687] = 32'h79baf248;
    ram_cell[     688] = 32'h918e5d9f;
    ram_cell[     689] = 32'hd4059e73;
    ram_cell[     690] = 32'ha45dbb63;
    ram_cell[     691] = 32'h563d2dac;
    ram_cell[     692] = 32'hcb35fe00;
    ram_cell[     693] = 32'h76d84119;
    ram_cell[     694] = 32'h682b5b88;
    ram_cell[     695] = 32'hd4f3f5e0;
    ram_cell[     696] = 32'hd58e1504;
    ram_cell[     697] = 32'h386993d3;
    ram_cell[     698] = 32'h70690248;
    ram_cell[     699] = 32'hb337fd12;
    ram_cell[     700] = 32'hde5de1b6;
    ram_cell[     701] = 32'h6dba8d0a;
    ram_cell[     702] = 32'h54214d77;
    ram_cell[     703] = 32'h6c114d85;
    ram_cell[     704] = 32'hcee51e3a;
    ram_cell[     705] = 32'hd7952a64;
    ram_cell[     706] = 32'he89c7290;
    ram_cell[     707] = 32'h8be0b23f;
    ram_cell[     708] = 32'h74acac5a;
    ram_cell[     709] = 32'h33da6ade;
    ram_cell[     710] = 32'h96737ba8;
    ram_cell[     711] = 32'h430e0373;
    ram_cell[     712] = 32'h53aaf7d9;
    ram_cell[     713] = 32'h682ff567;
    ram_cell[     714] = 32'h5f807792;
    ram_cell[     715] = 32'hf4bead65;
    ram_cell[     716] = 32'h0d4b1750;
    ram_cell[     717] = 32'h9d22970a;
    ram_cell[     718] = 32'hbe386450;
    ram_cell[     719] = 32'h3bde34c3;
    ram_cell[     720] = 32'hb5ad714d;
    ram_cell[     721] = 32'h75d848a4;
    ram_cell[     722] = 32'h9edbbe53;
    ram_cell[     723] = 32'hc1c12ed8;
    ram_cell[     724] = 32'h77a4a8ec;
    ram_cell[     725] = 32'hcaa6df15;
    ram_cell[     726] = 32'h4fb0256d;
    ram_cell[     727] = 32'h12c9197f;
    ram_cell[     728] = 32'h28e56e95;
    ram_cell[     729] = 32'h80726fbc;
    ram_cell[     730] = 32'hd14081f2;
    ram_cell[     731] = 32'he03949a8;
    ram_cell[     732] = 32'h4b04c86a;
    ram_cell[     733] = 32'hd4e64ef0;
    ram_cell[     734] = 32'h7fe2df7e;
    ram_cell[     735] = 32'habbd36aa;
    ram_cell[     736] = 32'h9c87fcb4;
    ram_cell[     737] = 32'h6ab55311;
    ram_cell[     738] = 32'h30746400;
    ram_cell[     739] = 32'h9379f308;
    ram_cell[     740] = 32'h0239faab;
    ram_cell[     741] = 32'hdd7c5274;
    ram_cell[     742] = 32'h1cda0413;
    ram_cell[     743] = 32'h9312532b;
    ram_cell[     744] = 32'h0a13d262;
    ram_cell[     745] = 32'h686e605f;
    ram_cell[     746] = 32'hb3a971e9;
    ram_cell[     747] = 32'h24d6aa01;
    ram_cell[     748] = 32'h8c2e7989;
    ram_cell[     749] = 32'h0b49fa62;
    ram_cell[     750] = 32'h1c7fac9b;
    ram_cell[     751] = 32'h5cd3662b;
    ram_cell[     752] = 32'h731eb7f6;
    ram_cell[     753] = 32'h6ee0a5c9;
    ram_cell[     754] = 32'h50f9da50;
    ram_cell[     755] = 32'hc264cda1;
    ram_cell[     756] = 32'hcae8f1de;
    ram_cell[     757] = 32'h52ecce7f;
    ram_cell[     758] = 32'ha691fa33;
    ram_cell[     759] = 32'h3bf62ebf;
    ram_cell[     760] = 32'h69f051d2;
    ram_cell[     761] = 32'h72ca5817;
    ram_cell[     762] = 32'hab82786f;
    ram_cell[     763] = 32'h638294f8;
    ram_cell[     764] = 32'he431778d;
    ram_cell[     765] = 32'h2ce34917;
    ram_cell[     766] = 32'hb10587e3;
    ram_cell[     767] = 32'h68ab9944;
end

endmodule

