
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'ha4898942;
    ram_cell[       1] = 32'h0;  // 32'h723ecc3a;
    ram_cell[       2] = 32'h0;  // 32'h1f078ce6;
    ram_cell[       3] = 32'h0;  // 32'ha478ddd7;
    ram_cell[       4] = 32'h0;  // 32'he255661a;
    ram_cell[       5] = 32'h0;  // 32'hf8176222;
    ram_cell[       6] = 32'h0;  // 32'h263ab724;
    ram_cell[       7] = 32'h0;  // 32'h815572e4;
    ram_cell[       8] = 32'h0;  // 32'h4568df74;
    ram_cell[       9] = 32'h0;  // 32'hef057ae9;
    ram_cell[      10] = 32'h0;  // 32'h4c577df6;
    ram_cell[      11] = 32'h0;  // 32'h64ad0423;
    ram_cell[      12] = 32'h0;  // 32'h93666dda;
    ram_cell[      13] = 32'h0;  // 32'hdf00d130;
    ram_cell[      14] = 32'h0;  // 32'h5668c07d;
    ram_cell[      15] = 32'h0;  // 32'h4776a5c2;
    ram_cell[      16] = 32'h0;  // 32'h93feb163;
    ram_cell[      17] = 32'h0;  // 32'h99ef0d1c;
    ram_cell[      18] = 32'h0;  // 32'hae1720bd;
    ram_cell[      19] = 32'h0;  // 32'h02cb7bb5;
    ram_cell[      20] = 32'h0;  // 32'haff74da1;
    ram_cell[      21] = 32'h0;  // 32'h5a26680d;
    ram_cell[      22] = 32'h0;  // 32'hcf3058e9;
    ram_cell[      23] = 32'h0;  // 32'h4a5293f6;
    ram_cell[      24] = 32'h0;  // 32'h14b26852;
    ram_cell[      25] = 32'h0;  // 32'h8a16a70d;
    ram_cell[      26] = 32'h0;  // 32'hfe3bccaf;
    ram_cell[      27] = 32'h0;  // 32'h2303358d;
    ram_cell[      28] = 32'h0;  // 32'h6e05604c;
    ram_cell[      29] = 32'h0;  // 32'hb1469b84;
    ram_cell[      30] = 32'h0;  // 32'hb6e91cc6;
    ram_cell[      31] = 32'h0;  // 32'h6b4694f8;
    ram_cell[      32] = 32'h0;  // 32'h676345ba;
    ram_cell[      33] = 32'h0;  // 32'h059b0335;
    ram_cell[      34] = 32'h0;  // 32'had1eeabd;
    ram_cell[      35] = 32'h0;  // 32'h9f13f100;
    ram_cell[      36] = 32'h0;  // 32'hc4ca22f3;
    ram_cell[      37] = 32'h0;  // 32'h82ef893f;
    ram_cell[      38] = 32'h0;  // 32'he293b312;
    ram_cell[      39] = 32'h0;  // 32'h5c8772d4;
    ram_cell[      40] = 32'h0;  // 32'h96cd29d7;
    ram_cell[      41] = 32'h0;  // 32'h3dc22a68;
    ram_cell[      42] = 32'h0;  // 32'hc78f186a;
    ram_cell[      43] = 32'h0;  // 32'h99f81e23;
    ram_cell[      44] = 32'h0;  // 32'h9e78286c;
    ram_cell[      45] = 32'h0;  // 32'h865e0efc;
    ram_cell[      46] = 32'h0;  // 32'h4e04228a;
    ram_cell[      47] = 32'h0;  // 32'h9f21efd3;
    ram_cell[      48] = 32'h0;  // 32'h3785a26b;
    ram_cell[      49] = 32'h0;  // 32'h405a0522;
    ram_cell[      50] = 32'h0;  // 32'h5df0b6e6;
    ram_cell[      51] = 32'h0;  // 32'ha5f9564d;
    ram_cell[      52] = 32'h0;  // 32'h64c1b5eb;
    ram_cell[      53] = 32'h0;  // 32'hc53d5244;
    ram_cell[      54] = 32'h0;  // 32'hd78fa1fe;
    ram_cell[      55] = 32'h0;  // 32'h8d1d646c;
    ram_cell[      56] = 32'h0;  // 32'h09cc1627;
    ram_cell[      57] = 32'h0;  // 32'hccbf7c36;
    ram_cell[      58] = 32'h0;  // 32'h9b12e2e5;
    ram_cell[      59] = 32'h0;  // 32'h4356690f;
    ram_cell[      60] = 32'h0;  // 32'h1a7c3dde;
    ram_cell[      61] = 32'h0;  // 32'h5cc4ce8d;
    ram_cell[      62] = 32'h0;  // 32'hfdc3db56;
    ram_cell[      63] = 32'h0;  // 32'haf6dff85;
    ram_cell[      64] = 32'h0;  // 32'h303ff1cc;
    ram_cell[      65] = 32'h0;  // 32'h583db0de;
    ram_cell[      66] = 32'h0;  // 32'h4c49c2a7;
    ram_cell[      67] = 32'h0;  // 32'hed610e04;
    ram_cell[      68] = 32'h0;  // 32'he6b2263a;
    ram_cell[      69] = 32'h0;  // 32'ha9d1f8b7;
    ram_cell[      70] = 32'h0;  // 32'hde0c9109;
    ram_cell[      71] = 32'h0;  // 32'hcc1a6163;
    ram_cell[      72] = 32'h0;  // 32'h06b9a265;
    ram_cell[      73] = 32'h0;  // 32'h36158a37;
    ram_cell[      74] = 32'h0;  // 32'heb3b0f1c;
    ram_cell[      75] = 32'h0;  // 32'ha224123f;
    ram_cell[      76] = 32'h0;  // 32'he387a426;
    ram_cell[      77] = 32'h0;  // 32'hd91a17ec;
    ram_cell[      78] = 32'h0;  // 32'h0299038b;
    ram_cell[      79] = 32'h0;  // 32'hcfc82a0f;
    ram_cell[      80] = 32'h0;  // 32'hfbf2e41d;
    ram_cell[      81] = 32'h0;  // 32'h3e036c79;
    ram_cell[      82] = 32'h0;  // 32'hc892b5ee;
    ram_cell[      83] = 32'h0;  // 32'h8cda4218;
    ram_cell[      84] = 32'h0;  // 32'h475beae1;
    ram_cell[      85] = 32'h0;  // 32'h4f96c3cc;
    ram_cell[      86] = 32'h0;  // 32'h01f20c92;
    ram_cell[      87] = 32'h0;  // 32'he233e44a;
    ram_cell[      88] = 32'h0;  // 32'h82c58ddf;
    ram_cell[      89] = 32'h0;  // 32'h4ddfe506;
    ram_cell[      90] = 32'h0;  // 32'hf7d90348;
    ram_cell[      91] = 32'h0;  // 32'hd48d1b6d;
    ram_cell[      92] = 32'h0;  // 32'hbd0cbc0a;
    ram_cell[      93] = 32'h0;  // 32'h3841a6c1;
    ram_cell[      94] = 32'h0;  // 32'ha18d57c7;
    ram_cell[      95] = 32'h0;  // 32'hb0ce396e;
    ram_cell[      96] = 32'h0;  // 32'hbc5ad20f;
    ram_cell[      97] = 32'h0;  // 32'h0c866fd4;
    ram_cell[      98] = 32'h0;  // 32'h6362dd5e;
    ram_cell[      99] = 32'h0;  // 32'h6e982553;
    ram_cell[     100] = 32'h0;  // 32'h485bf8a9;
    ram_cell[     101] = 32'h0;  // 32'hebcb63fa;
    ram_cell[     102] = 32'h0;  // 32'h3add499e;
    ram_cell[     103] = 32'h0;  // 32'h4e0dad6b;
    ram_cell[     104] = 32'h0;  // 32'haa9aa941;
    ram_cell[     105] = 32'h0;  // 32'h36483109;
    ram_cell[     106] = 32'h0;  // 32'hfd54942e;
    ram_cell[     107] = 32'h0;  // 32'h1d64f236;
    ram_cell[     108] = 32'h0;  // 32'h933c8adf;
    ram_cell[     109] = 32'h0;  // 32'h13938b8f;
    ram_cell[     110] = 32'h0;  // 32'ha6abe842;
    ram_cell[     111] = 32'h0;  // 32'hb7e95fd4;
    ram_cell[     112] = 32'h0;  // 32'h0f04e0f1;
    ram_cell[     113] = 32'h0;  // 32'he8f05cff;
    ram_cell[     114] = 32'h0;  // 32'ha7c1fa3d;
    ram_cell[     115] = 32'h0;  // 32'hbfd18843;
    ram_cell[     116] = 32'h0;  // 32'h6d891f6c;
    ram_cell[     117] = 32'h0;  // 32'hc3c3d14d;
    ram_cell[     118] = 32'h0;  // 32'h0ef2c5aa;
    ram_cell[     119] = 32'h0;  // 32'h0bb987d2;
    ram_cell[     120] = 32'h0;  // 32'h48728de9;
    ram_cell[     121] = 32'h0;  // 32'h70668044;
    ram_cell[     122] = 32'h0;  // 32'h95c7391b;
    ram_cell[     123] = 32'h0;  // 32'h8738d1e9;
    ram_cell[     124] = 32'h0;  // 32'h046ba99e;
    ram_cell[     125] = 32'h0;  // 32'h194a7b92;
    ram_cell[     126] = 32'h0;  // 32'h346624c6;
    ram_cell[     127] = 32'h0;  // 32'h7c51ddc1;
    ram_cell[     128] = 32'h0;  // 32'h19209bb8;
    ram_cell[     129] = 32'h0;  // 32'hf3ad46ac;
    ram_cell[     130] = 32'h0;  // 32'hed5622e6;
    ram_cell[     131] = 32'h0;  // 32'h2b6c2190;
    ram_cell[     132] = 32'h0;  // 32'h99840411;
    ram_cell[     133] = 32'h0;  // 32'h22aef36d;
    ram_cell[     134] = 32'h0;  // 32'h1dffc301;
    ram_cell[     135] = 32'h0;  // 32'h0b235a8b;
    ram_cell[     136] = 32'h0;  // 32'hcd936d81;
    ram_cell[     137] = 32'h0;  // 32'hc51736f9;
    ram_cell[     138] = 32'h0;  // 32'hc1848e2b;
    ram_cell[     139] = 32'h0;  // 32'h64333154;
    ram_cell[     140] = 32'h0;  // 32'h30d79765;
    ram_cell[     141] = 32'h0;  // 32'h6e8a1c7b;
    ram_cell[     142] = 32'h0;  // 32'h064f7b19;
    ram_cell[     143] = 32'h0;  // 32'h61cc9731;
    ram_cell[     144] = 32'h0;  // 32'h11b13e7c;
    ram_cell[     145] = 32'h0;  // 32'hc82db5c6;
    ram_cell[     146] = 32'h0;  // 32'h948733ac;
    ram_cell[     147] = 32'h0;  // 32'h4d0a31b4;
    ram_cell[     148] = 32'h0;  // 32'hf601611f;
    ram_cell[     149] = 32'h0;  // 32'hb4c2b2b2;
    ram_cell[     150] = 32'h0;  // 32'he7e915d2;
    ram_cell[     151] = 32'h0;  // 32'h6c4923c1;
    ram_cell[     152] = 32'h0;  // 32'hd44c57f1;
    ram_cell[     153] = 32'h0;  // 32'h792bd114;
    ram_cell[     154] = 32'h0;  // 32'h2ecd8950;
    ram_cell[     155] = 32'h0;  // 32'h0f3efa75;
    ram_cell[     156] = 32'h0;  // 32'he5a8ba66;
    ram_cell[     157] = 32'h0;  // 32'h7853dc46;
    ram_cell[     158] = 32'h0;  // 32'h393b3e74;
    ram_cell[     159] = 32'h0;  // 32'h5b66e1ba;
    ram_cell[     160] = 32'h0;  // 32'he9d42373;
    ram_cell[     161] = 32'h0;  // 32'h6ea1a414;
    ram_cell[     162] = 32'h0;  // 32'h8e3aa7e3;
    ram_cell[     163] = 32'h0;  // 32'h9e506be3;
    ram_cell[     164] = 32'h0;  // 32'h93847094;
    ram_cell[     165] = 32'h0;  // 32'hacec4a4d;
    ram_cell[     166] = 32'h0;  // 32'hc6a26829;
    ram_cell[     167] = 32'h0;  // 32'h70c15262;
    ram_cell[     168] = 32'h0;  // 32'hfb9f8e5d;
    ram_cell[     169] = 32'h0;  // 32'h0a625cf9;
    ram_cell[     170] = 32'h0;  // 32'h7e4be07e;
    ram_cell[     171] = 32'h0;  // 32'h50aae42d;
    ram_cell[     172] = 32'h0;  // 32'h41cca717;
    ram_cell[     173] = 32'h0;  // 32'hcc717169;
    ram_cell[     174] = 32'h0;  // 32'hac7cad26;
    ram_cell[     175] = 32'h0;  // 32'hc46950d9;
    ram_cell[     176] = 32'h0;  // 32'h8c181b60;
    ram_cell[     177] = 32'h0;  // 32'h84377fbb;
    ram_cell[     178] = 32'h0;  // 32'ha5851f4e;
    ram_cell[     179] = 32'h0;  // 32'h38d5b7b5;
    ram_cell[     180] = 32'h0;  // 32'hf65cb489;
    ram_cell[     181] = 32'h0;  // 32'hce593d7a;
    ram_cell[     182] = 32'h0;  // 32'h898bf0e3;
    ram_cell[     183] = 32'h0;  // 32'hf6191cbb;
    ram_cell[     184] = 32'h0;  // 32'h4789c5de;
    ram_cell[     185] = 32'h0;  // 32'h2df0d181;
    ram_cell[     186] = 32'h0;  // 32'h80f1db61;
    ram_cell[     187] = 32'h0;  // 32'h4f6f408d;
    ram_cell[     188] = 32'h0;  // 32'h560bba74;
    ram_cell[     189] = 32'h0;  // 32'h2a40854f;
    ram_cell[     190] = 32'h0;  // 32'h8517e752;
    ram_cell[     191] = 32'h0;  // 32'h1981e4e8;
    ram_cell[     192] = 32'h0;  // 32'he7371b71;
    ram_cell[     193] = 32'h0;  // 32'h9cff44b5;
    ram_cell[     194] = 32'h0;  // 32'hb229d6a4;
    ram_cell[     195] = 32'h0;  // 32'h76af2d6c;
    ram_cell[     196] = 32'h0;  // 32'h938c75d3;
    ram_cell[     197] = 32'h0;  // 32'h5cbc971a;
    ram_cell[     198] = 32'h0;  // 32'h075c0ad9;
    ram_cell[     199] = 32'h0;  // 32'h7d3c6ce9;
    ram_cell[     200] = 32'h0;  // 32'h4e0ea6a5;
    ram_cell[     201] = 32'h0;  // 32'h7d7eef12;
    ram_cell[     202] = 32'h0;  // 32'h21be1df1;
    ram_cell[     203] = 32'h0;  // 32'hf5bdb907;
    ram_cell[     204] = 32'h0;  // 32'hea3845f5;
    ram_cell[     205] = 32'h0;  // 32'h2392b9c1;
    ram_cell[     206] = 32'h0;  // 32'h12829241;
    ram_cell[     207] = 32'h0;  // 32'ha237e0b9;
    ram_cell[     208] = 32'h0;  // 32'h5bcccfd2;
    ram_cell[     209] = 32'h0;  // 32'hc662feab;
    ram_cell[     210] = 32'h0;  // 32'hb7436bbc;
    ram_cell[     211] = 32'h0;  // 32'h6a47de8b;
    ram_cell[     212] = 32'h0;  // 32'h6a994311;
    ram_cell[     213] = 32'h0;  // 32'hfdbb6ed1;
    ram_cell[     214] = 32'h0;  // 32'hf0f07ddd;
    ram_cell[     215] = 32'h0;  // 32'h67578446;
    ram_cell[     216] = 32'h0;  // 32'h12658e09;
    ram_cell[     217] = 32'h0;  // 32'h8ddb33b3;
    ram_cell[     218] = 32'h0;  // 32'hc87232e9;
    ram_cell[     219] = 32'h0;  // 32'hb595f5b4;
    ram_cell[     220] = 32'h0;  // 32'h381ff24b;
    ram_cell[     221] = 32'h0;  // 32'h0df9713e;
    ram_cell[     222] = 32'h0;  // 32'hdea10882;
    ram_cell[     223] = 32'h0;  // 32'h91865b99;
    ram_cell[     224] = 32'h0;  // 32'h97214f0f;
    ram_cell[     225] = 32'h0;  // 32'ha0d88ef2;
    ram_cell[     226] = 32'h0;  // 32'h1422cfec;
    ram_cell[     227] = 32'h0;  // 32'he33a7502;
    ram_cell[     228] = 32'h0;  // 32'he0094849;
    ram_cell[     229] = 32'h0;  // 32'haa0ffd41;
    ram_cell[     230] = 32'h0;  // 32'hc726e047;
    ram_cell[     231] = 32'h0;  // 32'h1e9a4c05;
    ram_cell[     232] = 32'h0;  // 32'hafc1d2d1;
    ram_cell[     233] = 32'h0;  // 32'h56d60f46;
    ram_cell[     234] = 32'h0;  // 32'h8081bcc3;
    ram_cell[     235] = 32'h0;  // 32'h015ebada;
    ram_cell[     236] = 32'h0;  // 32'hb4fd2431;
    ram_cell[     237] = 32'h0;  // 32'h4a9fa1e9;
    ram_cell[     238] = 32'h0;  // 32'he58df48d;
    ram_cell[     239] = 32'h0;  // 32'h1f46a0fe;
    ram_cell[     240] = 32'h0;  // 32'h36cd7a1f;
    ram_cell[     241] = 32'h0;  // 32'h4670bd4d;
    ram_cell[     242] = 32'h0;  // 32'h0085ff16;
    ram_cell[     243] = 32'h0;  // 32'hbfd5ab72;
    ram_cell[     244] = 32'h0;  // 32'h9f3b28b9;
    ram_cell[     245] = 32'h0;  // 32'h8da8630d;
    ram_cell[     246] = 32'h0;  // 32'h11dd7496;
    ram_cell[     247] = 32'h0;  // 32'h2c4c6816;
    ram_cell[     248] = 32'h0;  // 32'hca217fd6;
    ram_cell[     249] = 32'h0;  // 32'hcce3046b;
    ram_cell[     250] = 32'h0;  // 32'hd7ed0343;
    ram_cell[     251] = 32'h0;  // 32'h6f633d97;
    ram_cell[     252] = 32'h0;  // 32'ha5f35121;
    ram_cell[     253] = 32'h0;  // 32'h0f385488;
    ram_cell[     254] = 32'h0;  // 32'h661d7bbf;
    ram_cell[     255] = 32'h0;  // 32'h3e56b22d;
    // src matrix A
    ram_cell[     256] = 32'hf49940c5;
    ram_cell[     257] = 32'hab24676f;
    ram_cell[     258] = 32'h8e4a2e0a;
    ram_cell[     259] = 32'h725c3ebd;
    ram_cell[     260] = 32'h09e8fd9a;
    ram_cell[     261] = 32'h6e54ccd0;
    ram_cell[     262] = 32'hd667149a;
    ram_cell[     263] = 32'h83794803;
    ram_cell[     264] = 32'hfc2d82df;
    ram_cell[     265] = 32'h94d1e4c6;
    ram_cell[     266] = 32'hf2db8d26;
    ram_cell[     267] = 32'haf7d19a3;
    ram_cell[     268] = 32'h772c2b56;
    ram_cell[     269] = 32'h8232e107;
    ram_cell[     270] = 32'h009fdd2c;
    ram_cell[     271] = 32'h8464ac1b;
    ram_cell[     272] = 32'h3a127fd4;
    ram_cell[     273] = 32'hf2ff505d;
    ram_cell[     274] = 32'h164b2e12;
    ram_cell[     275] = 32'hdcbfd8dc;
    ram_cell[     276] = 32'h9ad7661e;
    ram_cell[     277] = 32'h9273fdab;
    ram_cell[     278] = 32'hee01522d;
    ram_cell[     279] = 32'hdc0af1ad;
    ram_cell[     280] = 32'h23f6a8c7;
    ram_cell[     281] = 32'hfba489a1;
    ram_cell[     282] = 32'h4837c666;
    ram_cell[     283] = 32'hc35ed59d;
    ram_cell[     284] = 32'h86c8cef0;
    ram_cell[     285] = 32'h1d59ee2e;
    ram_cell[     286] = 32'h02bc2ee7;
    ram_cell[     287] = 32'h80eb1c8b;
    ram_cell[     288] = 32'hda1854a4;
    ram_cell[     289] = 32'h5b475332;
    ram_cell[     290] = 32'hec81b24e;
    ram_cell[     291] = 32'haf6b4d04;
    ram_cell[     292] = 32'hf2640a38;
    ram_cell[     293] = 32'hcdd99839;
    ram_cell[     294] = 32'h63404e29;
    ram_cell[     295] = 32'h8ed413f0;
    ram_cell[     296] = 32'h875dfd70;
    ram_cell[     297] = 32'h0ce0bc78;
    ram_cell[     298] = 32'ha8ef3c09;
    ram_cell[     299] = 32'hf1a558e0;
    ram_cell[     300] = 32'h598fd394;
    ram_cell[     301] = 32'hf2d1cacf;
    ram_cell[     302] = 32'hb8ca1f8d;
    ram_cell[     303] = 32'h5eee0ed7;
    ram_cell[     304] = 32'h1cba8b6a;
    ram_cell[     305] = 32'h1da9855b;
    ram_cell[     306] = 32'hf99e623c;
    ram_cell[     307] = 32'h2d51023b;
    ram_cell[     308] = 32'hafc345e6;
    ram_cell[     309] = 32'h2eca4307;
    ram_cell[     310] = 32'h86ada128;
    ram_cell[     311] = 32'h00506b79;
    ram_cell[     312] = 32'h777d2b89;
    ram_cell[     313] = 32'h6d2d2cfc;
    ram_cell[     314] = 32'h9fbd29e9;
    ram_cell[     315] = 32'h7fbe8b54;
    ram_cell[     316] = 32'haa6c6dd3;
    ram_cell[     317] = 32'h2e9abe6f;
    ram_cell[     318] = 32'he8560021;
    ram_cell[     319] = 32'hf3cb0c97;
    ram_cell[     320] = 32'h3c1e38f9;
    ram_cell[     321] = 32'hebfe899e;
    ram_cell[     322] = 32'h1a3d2569;
    ram_cell[     323] = 32'he84d5f80;
    ram_cell[     324] = 32'h8bcb9e01;
    ram_cell[     325] = 32'h80e915c4;
    ram_cell[     326] = 32'h22fbcfc5;
    ram_cell[     327] = 32'h086228d1;
    ram_cell[     328] = 32'h08fbb00c;
    ram_cell[     329] = 32'h8a3aaeb3;
    ram_cell[     330] = 32'h7eea73a3;
    ram_cell[     331] = 32'h8aad4ae2;
    ram_cell[     332] = 32'h579f7e29;
    ram_cell[     333] = 32'h8f33c77a;
    ram_cell[     334] = 32'hefda99e6;
    ram_cell[     335] = 32'he16943f9;
    ram_cell[     336] = 32'hba5af72c;
    ram_cell[     337] = 32'h550b6689;
    ram_cell[     338] = 32'h43aeff69;
    ram_cell[     339] = 32'h86a44438;
    ram_cell[     340] = 32'h93bd657a;
    ram_cell[     341] = 32'he38b6d00;
    ram_cell[     342] = 32'h37d28151;
    ram_cell[     343] = 32'hdec1dc74;
    ram_cell[     344] = 32'h690cf7a2;
    ram_cell[     345] = 32'hde8b2544;
    ram_cell[     346] = 32'hc4e88d72;
    ram_cell[     347] = 32'h811100a1;
    ram_cell[     348] = 32'he00f497b;
    ram_cell[     349] = 32'h3611079f;
    ram_cell[     350] = 32'h9ef47142;
    ram_cell[     351] = 32'hc4aea010;
    ram_cell[     352] = 32'h6e491c78;
    ram_cell[     353] = 32'h895d8662;
    ram_cell[     354] = 32'h78a05add;
    ram_cell[     355] = 32'hc1bf3962;
    ram_cell[     356] = 32'h634f94eb;
    ram_cell[     357] = 32'h227e8620;
    ram_cell[     358] = 32'h1bded393;
    ram_cell[     359] = 32'h7319cbd5;
    ram_cell[     360] = 32'h63eacffb;
    ram_cell[     361] = 32'hc513211d;
    ram_cell[     362] = 32'h8dbc2709;
    ram_cell[     363] = 32'h4694f983;
    ram_cell[     364] = 32'h4dfacb52;
    ram_cell[     365] = 32'had7f567a;
    ram_cell[     366] = 32'hb2accce9;
    ram_cell[     367] = 32'h3d54869e;
    ram_cell[     368] = 32'h9f631ea0;
    ram_cell[     369] = 32'hed4b3363;
    ram_cell[     370] = 32'h1fd2ac71;
    ram_cell[     371] = 32'h7d0fb47c;
    ram_cell[     372] = 32'ha022ca9e;
    ram_cell[     373] = 32'h28614774;
    ram_cell[     374] = 32'hceeecc94;
    ram_cell[     375] = 32'he68c059d;
    ram_cell[     376] = 32'h93d1686d;
    ram_cell[     377] = 32'h37c58529;
    ram_cell[     378] = 32'h5be8004e;
    ram_cell[     379] = 32'h67cbaf14;
    ram_cell[     380] = 32'hdd3d39e8;
    ram_cell[     381] = 32'h11ec2004;
    ram_cell[     382] = 32'h9b6c6419;
    ram_cell[     383] = 32'h0a7d9291;
    ram_cell[     384] = 32'h71986744;
    ram_cell[     385] = 32'h62110e26;
    ram_cell[     386] = 32'h1f59afd2;
    ram_cell[     387] = 32'h442073b1;
    ram_cell[     388] = 32'h9009e21a;
    ram_cell[     389] = 32'h1a3588f1;
    ram_cell[     390] = 32'h52f6c3fd;
    ram_cell[     391] = 32'h68cc33b1;
    ram_cell[     392] = 32'h810379de;
    ram_cell[     393] = 32'h26157abb;
    ram_cell[     394] = 32'h21e0436e;
    ram_cell[     395] = 32'h8bad728f;
    ram_cell[     396] = 32'h24a5566f;
    ram_cell[     397] = 32'hfd1797db;
    ram_cell[     398] = 32'h96f02d05;
    ram_cell[     399] = 32'h6538eb94;
    ram_cell[     400] = 32'haa671542;
    ram_cell[     401] = 32'hb691c555;
    ram_cell[     402] = 32'h2ce7a679;
    ram_cell[     403] = 32'ha72655e8;
    ram_cell[     404] = 32'h6f753fa2;
    ram_cell[     405] = 32'h6894d8b4;
    ram_cell[     406] = 32'h7fb31cc8;
    ram_cell[     407] = 32'h11f6a1b0;
    ram_cell[     408] = 32'h36861dd7;
    ram_cell[     409] = 32'hb356c354;
    ram_cell[     410] = 32'h6befd6dc;
    ram_cell[     411] = 32'h3683f740;
    ram_cell[     412] = 32'h9d2a6104;
    ram_cell[     413] = 32'h2d90116c;
    ram_cell[     414] = 32'h4a1a660d;
    ram_cell[     415] = 32'hbf672c80;
    ram_cell[     416] = 32'h6a8bed63;
    ram_cell[     417] = 32'h721e475d;
    ram_cell[     418] = 32'h2bff186b;
    ram_cell[     419] = 32'h60203f07;
    ram_cell[     420] = 32'h346d1ffd;
    ram_cell[     421] = 32'h5d8adb1c;
    ram_cell[     422] = 32'hc12e3225;
    ram_cell[     423] = 32'hf7290543;
    ram_cell[     424] = 32'h36e3a061;
    ram_cell[     425] = 32'h6293a329;
    ram_cell[     426] = 32'h4ac44442;
    ram_cell[     427] = 32'hd32860c5;
    ram_cell[     428] = 32'h3f027d5e;
    ram_cell[     429] = 32'hf2e68ef2;
    ram_cell[     430] = 32'h8c5f838e;
    ram_cell[     431] = 32'hf18b951a;
    ram_cell[     432] = 32'h388a388e;
    ram_cell[     433] = 32'h604e4c0a;
    ram_cell[     434] = 32'he6c42daa;
    ram_cell[     435] = 32'h3407ff5f;
    ram_cell[     436] = 32'h5332d372;
    ram_cell[     437] = 32'h46e0f4ba;
    ram_cell[     438] = 32'h928f5b84;
    ram_cell[     439] = 32'h2db7afcd;
    ram_cell[     440] = 32'h3c9e007a;
    ram_cell[     441] = 32'h18e4e157;
    ram_cell[     442] = 32'h02afe9fb;
    ram_cell[     443] = 32'h37fb9972;
    ram_cell[     444] = 32'hb2415456;
    ram_cell[     445] = 32'h6431d18d;
    ram_cell[     446] = 32'hc73fed1a;
    ram_cell[     447] = 32'h5797b80b;
    ram_cell[     448] = 32'h632aabe4;
    ram_cell[     449] = 32'hbebba4e7;
    ram_cell[     450] = 32'h2e306ecc;
    ram_cell[     451] = 32'hdf705bc4;
    ram_cell[     452] = 32'hf1701895;
    ram_cell[     453] = 32'hcbc0b578;
    ram_cell[     454] = 32'h3aef2005;
    ram_cell[     455] = 32'h2cfe51c7;
    ram_cell[     456] = 32'h9e48e10b;
    ram_cell[     457] = 32'h7ed14a97;
    ram_cell[     458] = 32'h1bf39d2a;
    ram_cell[     459] = 32'hdb15a606;
    ram_cell[     460] = 32'hdca8d040;
    ram_cell[     461] = 32'hf3a2ffaa;
    ram_cell[     462] = 32'h528d6acf;
    ram_cell[     463] = 32'h6c6e558e;
    ram_cell[     464] = 32'h92c0134b;
    ram_cell[     465] = 32'h9b9e0224;
    ram_cell[     466] = 32'h310ba642;
    ram_cell[     467] = 32'hd143170a;
    ram_cell[     468] = 32'h8b2dd2f3;
    ram_cell[     469] = 32'h7c14631a;
    ram_cell[     470] = 32'ha70682f6;
    ram_cell[     471] = 32'h15ff91d9;
    ram_cell[     472] = 32'hb30379e3;
    ram_cell[     473] = 32'he579311d;
    ram_cell[     474] = 32'h3e560fd9;
    ram_cell[     475] = 32'hb5615ff1;
    ram_cell[     476] = 32'h2c0ebd39;
    ram_cell[     477] = 32'ha0286a0e;
    ram_cell[     478] = 32'h110ace04;
    ram_cell[     479] = 32'hd753a025;
    ram_cell[     480] = 32'h3cb27183;
    ram_cell[     481] = 32'hc0280ffe;
    ram_cell[     482] = 32'hd4b60f66;
    ram_cell[     483] = 32'h7933276a;
    ram_cell[     484] = 32'h415e7bbc;
    ram_cell[     485] = 32'hb1f20da1;
    ram_cell[     486] = 32'h27b85b70;
    ram_cell[     487] = 32'h4693bb3d;
    ram_cell[     488] = 32'h375e7695;
    ram_cell[     489] = 32'h9d0bed4e;
    ram_cell[     490] = 32'h9074711e;
    ram_cell[     491] = 32'he2f4a4db;
    ram_cell[     492] = 32'hda86d4ee;
    ram_cell[     493] = 32'hcc12b3cc;
    ram_cell[     494] = 32'h6c7f4e7e;
    ram_cell[     495] = 32'haa44d1ab;
    ram_cell[     496] = 32'hb5f72932;
    ram_cell[     497] = 32'hd08f99d8;
    ram_cell[     498] = 32'h9fc70456;
    ram_cell[     499] = 32'hef9fba38;
    ram_cell[     500] = 32'h02ead5c7;
    ram_cell[     501] = 32'hb824bd65;
    ram_cell[     502] = 32'h120ab082;
    ram_cell[     503] = 32'hc108b311;
    ram_cell[     504] = 32'h2e9c96d9;
    ram_cell[     505] = 32'h178a0dd8;
    ram_cell[     506] = 32'hb58f7261;
    ram_cell[     507] = 32'hd0039759;
    ram_cell[     508] = 32'h6d91efd2;
    ram_cell[     509] = 32'h2e412c79;
    ram_cell[     510] = 32'h08b909af;
    ram_cell[     511] = 32'he6e90753;
    // src matrix B
    ram_cell[     512] = 32'h8bc4cc9d;
    ram_cell[     513] = 32'h1c3306a7;
    ram_cell[     514] = 32'had5642a1;
    ram_cell[     515] = 32'h2842e2be;
    ram_cell[     516] = 32'h47611ddb;
    ram_cell[     517] = 32'h28ee193a;
    ram_cell[     518] = 32'hfde78dd9;
    ram_cell[     519] = 32'hcf3a6fb0;
    ram_cell[     520] = 32'h8aac3843;
    ram_cell[     521] = 32'h599a0439;
    ram_cell[     522] = 32'h9d821b64;
    ram_cell[     523] = 32'h0422fcb8;
    ram_cell[     524] = 32'hbfafd8f4;
    ram_cell[     525] = 32'he59975b6;
    ram_cell[     526] = 32'h96ecea65;
    ram_cell[     527] = 32'heffbc0dd;
    ram_cell[     528] = 32'h8ffa786c;
    ram_cell[     529] = 32'h1904e50c;
    ram_cell[     530] = 32'h7f03008a;
    ram_cell[     531] = 32'h00155903;
    ram_cell[     532] = 32'hc9f41328;
    ram_cell[     533] = 32'h4cb33d07;
    ram_cell[     534] = 32'h06e757d7;
    ram_cell[     535] = 32'h147597a8;
    ram_cell[     536] = 32'h27c100ea;
    ram_cell[     537] = 32'hfeb7d111;
    ram_cell[     538] = 32'h67a313d7;
    ram_cell[     539] = 32'h6f11987c;
    ram_cell[     540] = 32'hc76113fa;
    ram_cell[     541] = 32'h36fa1fa7;
    ram_cell[     542] = 32'he46fe778;
    ram_cell[     543] = 32'h9ab36c15;
    ram_cell[     544] = 32'h51d2f087;
    ram_cell[     545] = 32'h86a055f5;
    ram_cell[     546] = 32'heaffedf8;
    ram_cell[     547] = 32'h659ea59a;
    ram_cell[     548] = 32'h9c4c6f56;
    ram_cell[     549] = 32'h7fd6ad57;
    ram_cell[     550] = 32'h9ee0f04f;
    ram_cell[     551] = 32'h704df2e7;
    ram_cell[     552] = 32'h3dcd33fd;
    ram_cell[     553] = 32'h8d65425f;
    ram_cell[     554] = 32'h006244b7;
    ram_cell[     555] = 32'h4d40e0a8;
    ram_cell[     556] = 32'h6fe56ee0;
    ram_cell[     557] = 32'h82e64a02;
    ram_cell[     558] = 32'h6e20af41;
    ram_cell[     559] = 32'hebae9c60;
    ram_cell[     560] = 32'h50d194a6;
    ram_cell[     561] = 32'h26b26de0;
    ram_cell[     562] = 32'h52283fe4;
    ram_cell[     563] = 32'h1cc94d13;
    ram_cell[     564] = 32'h470524ba;
    ram_cell[     565] = 32'hbdb4efab;
    ram_cell[     566] = 32'h382d1e29;
    ram_cell[     567] = 32'hdcf4fe65;
    ram_cell[     568] = 32'h18a299d9;
    ram_cell[     569] = 32'h1473b174;
    ram_cell[     570] = 32'h11ed4dda;
    ram_cell[     571] = 32'he541a583;
    ram_cell[     572] = 32'h40f4da46;
    ram_cell[     573] = 32'h37ad3199;
    ram_cell[     574] = 32'hda1b5f8b;
    ram_cell[     575] = 32'hd190b70b;
    ram_cell[     576] = 32'h46ee1c33;
    ram_cell[     577] = 32'h2e3fcc97;
    ram_cell[     578] = 32'h43062986;
    ram_cell[     579] = 32'h6e66af1e;
    ram_cell[     580] = 32'h07d10ead;
    ram_cell[     581] = 32'hae4a2e0b;
    ram_cell[     582] = 32'h57a07235;
    ram_cell[     583] = 32'h202e187e;
    ram_cell[     584] = 32'h26e40a8e;
    ram_cell[     585] = 32'h8d472b93;
    ram_cell[     586] = 32'ha415e16e;
    ram_cell[     587] = 32'h037f9df1;
    ram_cell[     588] = 32'he7526a40;
    ram_cell[     589] = 32'hab9b814e;
    ram_cell[     590] = 32'ha73a6e77;
    ram_cell[     591] = 32'h9e6519d5;
    ram_cell[     592] = 32'hb10d49cc;
    ram_cell[     593] = 32'hcc1b8390;
    ram_cell[     594] = 32'h2ede4827;
    ram_cell[     595] = 32'he0c16a97;
    ram_cell[     596] = 32'h9dd88cbb;
    ram_cell[     597] = 32'h44686c6f;
    ram_cell[     598] = 32'hf6b41a08;
    ram_cell[     599] = 32'h5e8b8edf;
    ram_cell[     600] = 32'h05c6deb8;
    ram_cell[     601] = 32'h7d03c9eb;
    ram_cell[     602] = 32'hec9f1977;
    ram_cell[     603] = 32'h885f33c8;
    ram_cell[     604] = 32'h283993eb;
    ram_cell[     605] = 32'hc27a1b2c;
    ram_cell[     606] = 32'h880047f5;
    ram_cell[     607] = 32'h0c48faab;
    ram_cell[     608] = 32'h1b0cb9ec;
    ram_cell[     609] = 32'h758f2fd2;
    ram_cell[     610] = 32'h4bef1b63;
    ram_cell[     611] = 32'h9ea24a4a;
    ram_cell[     612] = 32'h14ad63b0;
    ram_cell[     613] = 32'h436a90e0;
    ram_cell[     614] = 32'h1945e0a6;
    ram_cell[     615] = 32'h68f9a929;
    ram_cell[     616] = 32'h963a741e;
    ram_cell[     617] = 32'h33f507ec;
    ram_cell[     618] = 32'h40578718;
    ram_cell[     619] = 32'h39410d59;
    ram_cell[     620] = 32'h0ed2e63b;
    ram_cell[     621] = 32'he8c14f7c;
    ram_cell[     622] = 32'h9fffe8d7;
    ram_cell[     623] = 32'h9ed838ed;
    ram_cell[     624] = 32'h200a53b9;
    ram_cell[     625] = 32'h7c4328e3;
    ram_cell[     626] = 32'h6586ad0a;
    ram_cell[     627] = 32'hae4b2613;
    ram_cell[     628] = 32'h5c20f216;
    ram_cell[     629] = 32'h5702f70a;
    ram_cell[     630] = 32'h2c8c8e56;
    ram_cell[     631] = 32'hd664fba0;
    ram_cell[     632] = 32'h68b93036;
    ram_cell[     633] = 32'h94dc9049;
    ram_cell[     634] = 32'hb2b763a7;
    ram_cell[     635] = 32'hc412b728;
    ram_cell[     636] = 32'h89ad36b8;
    ram_cell[     637] = 32'hdbe47f0e;
    ram_cell[     638] = 32'habdd47ae;
    ram_cell[     639] = 32'hc1aba0b5;
    ram_cell[     640] = 32'ha1058028;
    ram_cell[     641] = 32'hd5720da8;
    ram_cell[     642] = 32'heec9cfee;
    ram_cell[     643] = 32'h3b610d7e;
    ram_cell[     644] = 32'h5dff7ad9;
    ram_cell[     645] = 32'he6678c3f;
    ram_cell[     646] = 32'h115f3657;
    ram_cell[     647] = 32'h30c66ec6;
    ram_cell[     648] = 32'hb6477b9b;
    ram_cell[     649] = 32'h3dcc31b8;
    ram_cell[     650] = 32'hcf600b54;
    ram_cell[     651] = 32'h98245bb9;
    ram_cell[     652] = 32'h54ce0036;
    ram_cell[     653] = 32'hc5def620;
    ram_cell[     654] = 32'h0ea097a8;
    ram_cell[     655] = 32'hf744fd04;
    ram_cell[     656] = 32'h89f3004c;
    ram_cell[     657] = 32'hcbbb6824;
    ram_cell[     658] = 32'h777a147f;
    ram_cell[     659] = 32'hacd59d25;
    ram_cell[     660] = 32'h06a6a6ff;
    ram_cell[     661] = 32'h62b4b686;
    ram_cell[     662] = 32'he2461381;
    ram_cell[     663] = 32'h7b7b3ff0;
    ram_cell[     664] = 32'h2b5c2c57;
    ram_cell[     665] = 32'h13ae0bc1;
    ram_cell[     666] = 32'h398fe56d;
    ram_cell[     667] = 32'hb8a897e8;
    ram_cell[     668] = 32'hf79cfaae;
    ram_cell[     669] = 32'h5b56559f;
    ram_cell[     670] = 32'h7ac5af80;
    ram_cell[     671] = 32'hbaca15f6;
    ram_cell[     672] = 32'h86f975e4;
    ram_cell[     673] = 32'h2362b93a;
    ram_cell[     674] = 32'hec4d43bc;
    ram_cell[     675] = 32'h158ef1df;
    ram_cell[     676] = 32'he838022a;
    ram_cell[     677] = 32'h66cdfc90;
    ram_cell[     678] = 32'ha040a077;
    ram_cell[     679] = 32'hd36c2bb6;
    ram_cell[     680] = 32'hb1961ad5;
    ram_cell[     681] = 32'h9c837fca;
    ram_cell[     682] = 32'h2d1b277b;
    ram_cell[     683] = 32'ha3b88454;
    ram_cell[     684] = 32'h8b3d5114;
    ram_cell[     685] = 32'he4a2289f;
    ram_cell[     686] = 32'h1f33168f;
    ram_cell[     687] = 32'h637e0547;
    ram_cell[     688] = 32'he53bc4db;
    ram_cell[     689] = 32'he7d7802c;
    ram_cell[     690] = 32'hd9f1c8ce;
    ram_cell[     691] = 32'he4f209b1;
    ram_cell[     692] = 32'h7c56eece;
    ram_cell[     693] = 32'h5f7b238e;
    ram_cell[     694] = 32'hc7021b42;
    ram_cell[     695] = 32'h1c45c625;
    ram_cell[     696] = 32'h221df3e0;
    ram_cell[     697] = 32'he7553201;
    ram_cell[     698] = 32'he6227f96;
    ram_cell[     699] = 32'h7a427df7;
    ram_cell[     700] = 32'hae980528;
    ram_cell[     701] = 32'h75cbb140;
    ram_cell[     702] = 32'hdc35d4b5;
    ram_cell[     703] = 32'h5e570f3f;
    ram_cell[     704] = 32'hc6e443ee;
    ram_cell[     705] = 32'he00cb970;
    ram_cell[     706] = 32'h9eff9a4e;
    ram_cell[     707] = 32'h7e7c1b48;
    ram_cell[     708] = 32'hb1e4c0cf;
    ram_cell[     709] = 32'h29271268;
    ram_cell[     710] = 32'h493d5e37;
    ram_cell[     711] = 32'hb6353162;
    ram_cell[     712] = 32'heb40edf2;
    ram_cell[     713] = 32'hcfd2f1ea;
    ram_cell[     714] = 32'h30990aad;
    ram_cell[     715] = 32'h37ee2eb9;
    ram_cell[     716] = 32'h492c810b;
    ram_cell[     717] = 32'hbc1fd121;
    ram_cell[     718] = 32'h61395994;
    ram_cell[     719] = 32'h56f6afec;
    ram_cell[     720] = 32'hb655a4b5;
    ram_cell[     721] = 32'h8e16e1f2;
    ram_cell[     722] = 32'h889c3deb;
    ram_cell[     723] = 32'ha2bb0068;
    ram_cell[     724] = 32'h1354e60c;
    ram_cell[     725] = 32'hd633e3a2;
    ram_cell[     726] = 32'h649b5f3d;
    ram_cell[     727] = 32'h935b746d;
    ram_cell[     728] = 32'h38141250;
    ram_cell[     729] = 32'h106ff045;
    ram_cell[     730] = 32'h5a524b5d;
    ram_cell[     731] = 32'hc72c801a;
    ram_cell[     732] = 32'hd3191a3a;
    ram_cell[     733] = 32'hd76e044d;
    ram_cell[     734] = 32'h0ad57b58;
    ram_cell[     735] = 32'h0b7e8155;
    ram_cell[     736] = 32'hab3c6d8b;
    ram_cell[     737] = 32'h206fc033;
    ram_cell[     738] = 32'hd499341c;
    ram_cell[     739] = 32'h77eb1ead;
    ram_cell[     740] = 32'hc37f05e8;
    ram_cell[     741] = 32'hbdda0471;
    ram_cell[     742] = 32'h667b3df1;
    ram_cell[     743] = 32'hf57a260e;
    ram_cell[     744] = 32'hd423ef59;
    ram_cell[     745] = 32'hfc1345e4;
    ram_cell[     746] = 32'hefc06cd4;
    ram_cell[     747] = 32'haa30a324;
    ram_cell[     748] = 32'h7e5f2f1a;
    ram_cell[     749] = 32'h1f45b92f;
    ram_cell[     750] = 32'h99738f8d;
    ram_cell[     751] = 32'h87ae0111;
    ram_cell[     752] = 32'h44249a4a;
    ram_cell[     753] = 32'h5c287b32;
    ram_cell[     754] = 32'h1b93993a;
    ram_cell[     755] = 32'hd7484009;
    ram_cell[     756] = 32'he423f0fc;
    ram_cell[     757] = 32'h5dd4c07b;
    ram_cell[     758] = 32'h0269ed5f;
    ram_cell[     759] = 32'hf7f17987;
    ram_cell[     760] = 32'h6b0896f7;
    ram_cell[     761] = 32'ha5aabd8c;
    ram_cell[     762] = 32'hb93db2b7;
    ram_cell[     763] = 32'hb9cccdd4;
    ram_cell[     764] = 32'hdb5e05e6;
    ram_cell[     765] = 32'h3cbe1109;
    ram_cell[     766] = 32'haa4ff9c2;
    ram_cell[     767] = 32'hfd40cf9a;
end

endmodule

